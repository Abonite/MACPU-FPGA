module ddr3 (
);
    
endmodule