module mba (
    
);