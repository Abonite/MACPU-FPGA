`define	NOP         16'h0
`define	MOV_AR      16'h1
`define	MOV_RR      16'h2
`define	MOV_RA      16'h3
`define	LOAD        16'h4
`define	ADD_RR      16'h10
`define	ADD_RI      16'h110
`define	SUB_RR      16'h11
`define	SUB_RI      16'h111
`define	AND_RR      16'h12
`define	AND_RI      16'h112
`define	OR_RR       16'h13
`define	OR_RI       16'h113
`define	NOT_RR      16'h14
`define	NOT_RI      16'h114
`define	XOR_RR      16'h15
`define	XOR_RI      16'h115
`define	RAND_R      16'h16
`define	RAND_I      16'h116
`define	ROR_R       16'h17
`define	ROR_I       16'h117
`define	RXOR_R      16'h18
`define	RXOR_I      16'h118
`define	LSL_R       16'h19
`define	LSL_I       16'h119
`define	LSR_R       16'h1a
`define	LSR_I       16'h11a
`define	ASL_R       16'h1b
`define	ASL_I       16'h11b
`define	ASR_R       16'h1c
`define	ASR_I       16'h11c
`define	CSL_R       16'h1d
`define	CSL_I       16'h11d
`define	CSR_R       16'h1e
`define	CSR_I       16'h11e
`define	INC         16'h1f
`define	DEC         16'h20
`define	JMP         16'h40
`define	PUSH        16'h50
`define	POP         16'h51
`define	INT         16'h80
`define	SAVEPC      16'h81
`define	RECOPC      16'h82
