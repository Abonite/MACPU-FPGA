`define NOP         16'h0
`define MOV_AR      16'h1
`define MOV_RR      16'h2
`define MOV_RA      16'h3
`define LOAD        16'h4
`define ADD         16'h100
`define SUB         16'h101
`define AND         16'h102
`define OR          16'h103
`define NOT         16'h104
`define XOR         16'h105
`define RAND        16'h106
`define ROR         16'h107
`define RXOR        16'h108
`define LSL         16'h109
`define LSR         16'h10A
`define ASL         16'h10B
`define ASR         16'h10C
`define CSL         16'h10D
`define CSR         16'h10E
`define INC         16'h110
`define DEC         16'h111
`define JMP         16'h200
`define JMP         16'h200
`define PUSH        16'h400
`define POP         16'h401
`define INT         16'h8000
